<svg xmlns="http://www.w3.org/2000/svg" width="55" height="55" viewBox="0 0 55 55">
    <g fill="#FFF" fill-rule="evenodd">
        <path d="M2.316 52.464l.416-37.8h49.296l-.416 37.8H2.316zm49.847-50.11l-.11 9.955H2.88V2.354h49.283zm2.307-1.266c-.003-.046-.005-.094-.014-.14-.008-.039-.02-.075-.033-.112-.01-.036-.018-.073-.032-.109-.016-.04-.04-.077-.06-.116-.016-.029-.028-.059-.046-.085-.028-.045-.063-.084-.098-.123-.014-.018-.026-.038-.041-.054l-.002-.002A1.189 1.189 0 0 0 53.97.2c-.01-.008-.022-.012-.034-.019a1.119 1.119 0 0 0-.164-.091c-.02-.009-.041-.013-.063-.02-.05-.018-.1-.036-.153-.047a1.11 1.11 0 0 0-.23-.024H1.729c-.079 0-.156.008-.23.024-.02.004-.039.013-.06.018-.052.014-.106.029-.157.05-.017.008-.033.019-.05.027-.05.025-.1.05-.145.081-.018.012-.033.028-.05.042-.042.032-.083.063-.12.1-.018.02-.032.042-.05.061C.837.44.803.476.777.516.758.542.745.572.73.6.709.637.686.674.67.714.656.747.648.784.637.818.626.856.61.893.602.934c-.007.035-.008.072-.012.108-.004.04-.013.08-.013.122L0 53.627c-.003.315.117.618.333.841.216.224.512.35.819.35H52.75c.632 0 1.145-.52 1.152-1.164l.435-39.615c.087-.165.14-.352.14-.553V1.177c0-.03-.006-.059-.008-.089z"/>
        <path d="M7.534 6.55a1.064 1.064 0 0 1 1.532 0c.205.209.317.486.317.781 0 .296-.112.574-.317.782a1.09 1.09 0 0 1-1.532 0 1.105 1.105 0 0 1-.317-.782c0-.295.112-.572.317-.782m.767 4.241c.866 0 1.733-.336 2.393-1.011.64-.654.992-1.523.992-2.448 0-.924-.352-1.793-.992-2.446a3.335 3.335 0 0 0-4.788 0 3.476 3.476 0 0 0-.992 2.446c0 .925.353 1.794.992 2.447a3.334 3.334 0 0 0 2.395 1.012M15.281 6.55a1.063 1.063 0 0 1 1.532 0c.205.209.317.486.317.781 0 .296-.112.574-.317.782a1.09 1.09 0 0 1-1.532 0 1.105 1.105 0 0 1-.317-.782c0-.295.112-.572.317-.782m.766 4.241c.867 0 1.735-.336 2.394-1.012.64-.653.992-1.522.992-2.447 0-.924-.352-1.793-.992-2.446a3.336 3.336 0 0 0-4.788 0 3.476 3.476 0 0 0-.992 2.446c0 .925.352 1.794.992 2.447a3.333 3.333 0 0 0 2.394 1.012M23.028 6.55a1.064 1.064 0 0 1 1.532 0c.205.209.317.486.317.781 0 .296-.112.574-.317.782a1.09 1.09 0 0 1-1.532 0 1.105 1.105 0 0 1-.317-.782c0-.295.112-.572.317-.782m.766 4.241c.867 0 1.734-.336 2.394-1.011.64-.654.992-1.523.992-2.448 0-.924-.352-1.793-.992-2.446a3.335 3.335 0 0 0-4.788 0 3.476 3.476 0 0 0-.992 2.446c0 .925.352 1.794.992 2.447a3.334 3.334 0 0 0 2.394 1.012M37.658 35.416a1.144 1.144 0 0 0-.07.08l-2.528 2.583-1.787-1.827 2.598-2.655a1.196 1.196 0 0 0-.003-1.667l-2.595-2.653 1.787-1.827 5.196 5.31-2.598 2.656zm-1.784-10.463a1.14 1.14 0 0 0-.814-.344 1.14 1.14 0 0 0-.814.344l-3.416 3.491c-.216.221-.337.52-.337.833 0 .312.12.611.337.832l2.598 2.655-2.598 2.656a1.19 1.19 0 0 0-.337.832c0 .312.12.612.337.832l3.416 3.49a1.135 1.135 0 0 0 1.628 0l3.415-3.49c.025-.025.049-.051.07-.079l3.339-3.412c.45-.46.45-1.204 0-1.664l-6.824-6.976zM19.42 38.078l-2.548-2.6a1.268 1.268 0 0 0-.053-.059l-2.596-2.652 2.599-2.655c.023-.024.046-.048.067-.073l2.53-2.589 1.787 1.827-2.598 2.655c-.45.46-.446 1.208.003 1.667l2.595 2.653-1.787 1.826zm4.23-2.659l-2.599-2.654 2.598-2.656c.45-.46.45-1.204 0-1.664l-3.415-3.492a1.168 1.168 0 0 0-1.629 0l-3.414 3.492c-.024.023-.046.049-.067.074l-3.343 3.416a1.191 1.191 0 0 0 0 1.664l6.824 6.976c.217.22.51.345.815.345.305 0 .598-.124.814-.345l3.415-3.492c.45-.46.45-1.204 0-1.664zM29.01 19.681c-.625-.108-1.22.328-1.324.97l-3.854 23.844c-.104.641.321 1.247.948 1.353a1.158 1.158 0 0 0 1.324-.97l3.854-23.844a1.173 1.173 0 0 0-.948-1.353"/>
    </g>
</svg>
